../CPU/phymem.vhd