../CPU/alu.vhd