../CPU/decode.vhd