../CPU/cpu.vhd